library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity pattern_generator is
    Port (
        -- inputs
        clk                 : in std_logic;
        reset               : in std_logic;
        FIFO_full           : in std_logic;
        FIFO_wr_busy        : in std_logic;
        --VGA_VSYNC           : in std_logic_vector(11 downto 0);
        
        -- outputs
        -- signals handling color intensity
        gen_pixel             : out std_logic_vector(11 downto 0);
        FIFO_wr_en            : out std_logic
        -- signals handling frame printing
        --requested_pixel     : out std_logic_vector(11 downto 0); -- get the requested pixel from a frame buffer
    );
end pattern_generator;

architecture Behavioral of pattern_generator is

    signal cmp_end_line             : std_logic;
    signal cmp_end_frame            : std_logic;
    
    -- counters signal
    -- cols counter
    signal col_cnt                  : unsigned(9 downto 0);
    signal row_cnt                  : unsigned(9 downto 0);
    
    -- LUT signals for 'chess board' test pattern
    signal square                   : std_logic := '1';
    signal change_square            : unsigned(9 downto 0);
    signal square1                  : std_logic := '1';
    signal square2                  : std_logic := '0';
    signal invert_row               : std_logic := '0';
    constant square_width           : positive := 40;
    
begin

    process(clk, reset)
    begin
        if (reset = '1') then
            col_cnt <= to_unsigned(0, 10);
            row_cnt <= to_unsigned(0, 10);

        elsif (rising_edge(clk)) then
            -- cols counter logic
            if (cmp_end_line = '1') then
                col_cnt <= to_unsigned(0, 10);
            -- increment the cols at each clock cycle
            -- if the FIFO is not full or not busy
            elsif (fifo_full = '0') then
                col_cnt <= col_cnt + 1;
            end if;

            -- rows counter logic
            if (cmp_end_frame = '1') then
                row_cnt <= to_unsigned(0, 10);
            -- increment the rows when col_cnt = 639
            elsif (cmp_end_line = '1') then
                row_cnt <= row_cnt + 1;
            end if;

        end if;
    end process;

    -- combinatory logic

    --- LUT begining
    --- RGB test pattern
    gen_pixel <= x"000" when col_cnt < 320
        else x"FFF";
    --- LUT end

    --- LUT begining
    --- RGB test pattern
--    gen_pixel <= x"F00" when col_cnt < 160
--        else x"0F0" when col_cnt >= 160 and col_cnt < 320
--        else x"00F" when col_cnt >= 320 and col_cnt < 480
--        else x"FFF" when col_cnt >= 480 and col_cnt < 640;
    --- LUT end
    
    --- LUT begining
    --- RGB test pattern
--    gen_pixel <= (others => square);
    
    -- alternate square on row each 40 cols
--    change_square <= col_cnt mod square_width; -- square_width = 40
--    square <= not square when change_square = 0 else square;
    
    -- alternate square on col each 40 rows
--    invert_row <= '1' when row_cnt mod square_width = 0 else '0';
    
--    process(col_cnt, row_cnt)
--    begin
--        -- alternate square on row each 40 cols
--        if (col_cnt mod square_width = 0) then
--            square <= not square;
--        end if;
        
--        -- alternate square on col each 40 rows
--        if (row_cnt mod square_width = 0) then
--            invert_row <= not invert_row;
--        end if;
--    end process;
    
--    gen_pixel <= (others => square);-- when invert_row = '0' else (others => not square);
    
    --- LUT end
    
    cmp_end_line <= '1' when col_cnt = 639 else '0';
    cmp_end_frame <= '1' when row_cnt = 479 and col_cnt = 639 else '0';
    
    -- 
    FIFO_wr_en <= '1' when (col_cnt < 640 and row_cnt < 480) and (FIFO_full = '0') else '0';


end Behavioral;
